module backend

import v2.ast
import strings

pub struct CleanCGen {
	file ast.File
mut:
	sb        strings.Builder
	indent    int
	fn_types  map[string]string
	var_types map[string]string
}

pub fn CleanCGen.new(file ast.File) &CleanCGen {
	mut g := &CleanCGen{
		file:      file
		sb:        strings.new_builder(4096)
		fn_types:  map[string]string{}
		var_types: map[string]string{}
	}
	// Pass 0: Register function return types
	for stmt in file.stmts {
		if stmt is ast.FnDecl {
			mut ret := 'void'
			if stmt.typ.str() != 'void' && stmt.typ.str() != '' {
				ret = g.type_to_c(stmt.typ)
			}
			g.fn_types[stmt.name] = ret
		}
	}
	return g
}

pub fn (mut g CleanCGen) gen() string {
	g.sb.writeln('// Generated by V Clean C Backend')
	g.sb.writeln('#include <stdio.h>')
	g.sb.writeln('#include <stdlib.h>')
	g.sb.writeln('#include <stdbool.h>')
	g.sb.writeln('#include <stdint.h>')
	g.sb.writeln('')

	g.sb.writeln('typedef struct { char* str; int len; } string;')
	g.sb.writeln('')

	// 1. Struct Declarations (Typedefs)
	for stmt in g.file.stmts {
		if stmt is ast.StructDecl {
			g.sb.writeln('typedef struct ${stmt.name} ${stmt.name};')
		}
	}
	g.sb.writeln('')

	// 2. Struct Definitions
	for stmt in g.file.stmts {
		if stmt is ast.StructDecl {
			g.gen_struct_decl(stmt)
			g.sb.writeln('')
		}
	}

	// 3. Globals
	for stmt in g.file.stmts {
		if stmt is ast.GlobalDecl {
			g.gen_global_decl(stmt)
			g.sb.writeln('')
		}
	}

	// 4. Function Prototypes
	for stmt in g.file.stmts {
		if stmt is ast.FnDecl {
			g.gen_fn_head(stmt)
			g.sb.writeln(';')
		}
	}
	g.sb.writeln('')

	// 5. Functions
	for stmt in g.file.stmts {
		if stmt is ast.FnDecl {
			g.gen_fn_decl(stmt)
			g.sb.writeln('')
		}
	}

	return g.sb.str()
}

fn (mut g CleanCGen) type_to_c(t ast.Type) string {
	s := t.str()
	if s == 'string' {
		return 'string'
	}
	return s
}

fn (mut g CleanCGen) infer_type(node ast.Expr) string {
	match node {
		ast.BasicLiteral {
			if node.kind == .number {
				return 'int'
			}
			if node.kind in [.key_true, .key_false] {
				return 'bool'
			}
		}
		ast.StringLiteral {
			if node.value.starts_with("c'") {
				return 'char*'
			}
			return 'string'
		}
		ast.InitExpr {
			return node.typ.str()
		}
		ast.CallExpr {
			mut name := ''
			if node.lhs is ast.Ident {
				name = node.lhs.name
			} else if node.lhs is ast.SelectorExpr {
				name = node.lhs.rhs.name
			}

			if t := g.fn_types[name] {
				return t
			}
			// C builtins defaults
			if name in ['printf', 'puts', 'putchar'] {
				return 'int'
			}
			return 'int'
		}
		ast.Ident {
			if t := g.var_types[node.name] {
				return t
			}
			return 'int'
		}
		ast.ParenExpr {
			return g.infer_type(node.expr)
		}
		ast.InfixExpr {
			return g.infer_type(node.lhs)
		}
		else {
			return 'int'
		}
	}
	return ''
}

fn (mut g CleanCGen) gen_struct_decl(node ast.StructDecl) {
	g.sb.writeln('struct ${node.name} {')
	for field in node.fields {
		g.write_indent()
		g.sb.write_string('\t')
		t := 'field_type' // g.type_to_c(field.typ)
		g.sb.writeln('${t} ${field.name};')
	}
	g.sb.writeln('};')
}

fn (mut g CleanCGen) gen_global_decl(node ast.GlobalDecl) {
	for field in node.fields {
		t := 'field_type' // g.type_to_c(field.typ)
		g.sb.writeln('${t} ${field.name};')
	}
}

fn (mut g CleanCGen) gen_fn_head(node ast.FnDecl) {
	mut ret := 'void'
	if node.typ.str() != 'void' && node.typ.str() != '' {
		ret = g.type_to_c(node.typ)
	}
	if node.name == 'main' {
		ret = 'int'
	}
	g.sb.write_string('${ret} ${node.name}(')
	for i, param in node.typ.params {
		if i > 0 {
			g.sb.write_string(', ')
		}
		t := 'TYPE' // g.type_to_c(param.typ)
		g.sb.write_string('${t} ${param.name}')
	}
	g.sb.write_string(')')
}

fn (mut g CleanCGen) gen_fn_decl(node ast.FnDecl) {
	g.var_types = map[string]string{}
	// Register params
	for param in node.typ.params {
		g.var_types[param.name] = 'TYPE' // g.type_to_c(param.typ)
	}

	g.gen_fn_head(node)
	g.sb.writeln(' {')
	g.indent++
	g.gen_stmts(node.stmts)

	if node.name == 'main' {
		g.write_indent()
		g.sb.writeln('return 0;')
	}
	g.indent--
	g.sb.writeln('}')
}

fn (mut g CleanCGen) gen_stmts(stmts []ast.Stmt) {
	for s in stmts {
		g.gen_stmt(s)
	}
}

fn (mut g CleanCGen) gen_stmt(node ast.Stmt) {
	match node {
		ast.AssignStmt {
			g.write_indent()
			lhs := node.lhs[0]
			rhs := node.rhs[0]
			if node.op == .decl_assign {
				// var decl
				mut name := ''
				if lhs is ast.Ident {
					name = lhs.name
				}
				typ := g.infer_type(rhs)
				g.var_types[name] = typ
				g.sb.write_string('${typ} ${name} = ')
				g.gen_expr(rhs)
				g.sb.writeln(';')
			} else {
				// assignment
				g.gen_expr(lhs)
				op_str := match node.op {
					.assign { '=' }
					.plus_assign { '+=' }
					.minus_assign { '-=' }
					else { '=' }
				}
				g.sb.write_string(' ${op_str} ')
				g.gen_expr(rhs)
				g.sb.writeln(';')
			}
		}
		ast.ExprStmt {
			g.write_indent()
			g.gen_expr(node.expr)
			g.sb.writeln(';')
		}
		ast.ReturnStmt {
			g.write_indent()
			g.sb.write_string('return')
			if node.exprs.len > 0 {
				g.sb.write_string(' ')
				g.gen_expr(node.exprs[0])
			}
			g.sb.writeln(';')
		}
		ast.BlockStmt {
			g.write_indent()
			g.sb.writeln('{')
			g.indent++
			g.gen_stmts(node.stmts)
			g.indent--
			g.write_indent()
			g.sb.writeln('}')
		}
		ast.ForStmt {
			g.write_indent()
			if node.init is ast.EmptyStmt && node.cond is ast.EmptyExpr
				&& node.post is ast.EmptyStmt {
				g.sb.writeln('while (1) {')
			} else if node.init is ast.EmptyStmt && node.post is ast.EmptyStmt {
				g.sb.write_string('while (')
				g.gen_expr(node.cond)
				g.sb.writeln(') {')
			} else {
				g.sb.write_string('for (')
				if node.init !is ast.EmptyStmt {
					g.gen_stmt_inline(node.init)
				}
				g.sb.write_string('; ')
				if node.cond !is ast.EmptyExpr {
					g.gen_expr(node.cond)
				}
				g.sb.write_string('; ')
				if node.post !is ast.EmptyStmt {
					g.gen_stmt_inline(node.post)
				}
				g.sb.writeln(') {')
			}
			g.indent++
			g.gen_stmts(node.stmts)
			g.indent--
			g.write_indent()
			g.sb.writeln('}')
		}
		ast.FlowControlStmt {
			g.write_indent()
			if node.op == .key_break {
				g.sb.writeln('break;')
			} else {
				g.sb.writeln('continue;')
			}
		}
		else {
			g.sb.writeln('// Unhandled stmt: ${node.type_name()}')
		}
	}
}

fn (mut g CleanCGen) gen_stmt_inline(node ast.Stmt) {
	match node {
		ast.AssignStmt {
			lhs := node.lhs[0]
			rhs := node.rhs[0]
			if node.op == .decl_assign {
				mut name := ''
				if lhs is ast.Ident {
					name = lhs.name
				}
				t := g.infer_type(rhs)
				g.var_types[name] = t
				g.sb.write_string('${t} ${name} = ')
				g.gen_expr(rhs)
			} else {
				g.gen_expr(lhs)
				op := match node.op {
					.assign { '=' }
					.plus_assign { '+=' }
					.minus_assign { '-=' }
					else { '=' }
				}
				g.sb.write_string(' ${op} ')
				g.gen_expr(rhs)
			}
		}
		ast.ExprStmt {
			g.gen_expr(node.expr)
		}
		else {}
	}
}

fn (mut g CleanCGen) gen_expr(node ast.Expr) {
	match node {
		ast.BasicLiteral {
			if node.kind == .key_true {
				g.sb.write_string('true')
			} else if node.kind == .key_false {
				g.sb.write_string('false')
			} else {
				g.sb.write_string(node.value)
			}
		}
		ast.StringLiteral {
			if node.value.starts_with("c'") {
				val := node.value.trim("c'").trim("'")
				g.sb.write_string('"${val}"')
			} else {
				val := node.value.trim("'").trim('"')
				g.sb.write_string('(string){"${val}", ${val.len}}')
			}
		}
		ast.Ident {
			g.sb.write_string(node.name)
		}
		ast.IfExpr {
			// Statement IF
			g.write_indent()
			g.sb.write_string('if (')
			g.gen_expr(node.cond)
			g.sb.writeln(') {')
			g.indent++
			g.gen_stmts(node.stmts)
			g.indent--
			g.write_indent()
			g.sb.writeln('}')
			/*
			if node.else_stmts.len > 0 || node.else_expr !is ast.EmptyExpr {
				g.write_indent()
				g.sb.write_string('else ')
				if node.else_expr !is ast.EmptyExpr {
					// Inline else if
					// Cast expr to stmt implicitly by handling it inline
					// We need to print it without newline if possible?
					// Actually gen_stmt prints indent.
					// We hack it:
					// Treat else_expr (which is IfExpr) as a construct
					// We cannot call gen_stmt because it adds indent and newline.
					// Recursively handle the if part.
					// But for simplicity, let's just open a block or handle it.
					// Since we can't easily recurse without indent, block is safer.
					g.sb.writeln('{')
					g.indent++
					g.gen_stmt(ast.Stmt(node.else_expr))
					g.indent--
					g.write_indent()
					g.sb.writeln('}')
				} else {
					g.sb.writeln('{')
					g.indent++
					g.gen_stmts(node.else_stmts)
					g.indent--
					g.write_indent()
					g.sb.writeln('}')
				}
			}
			*/
		}
		ast.MatchExpr {
			g.write_indent()
			g.sb.write_string('switch (')
			g.gen_expr(node.expr)
			g.sb.writeln(') {')
			for branch in node.branches {
				if branch.cond.len == 0 {
					g.write_indent()
					g.sb.writeln('default:')
				} else {
					for c in branch.cond {
						g.write_indent()
						g.sb.write_string('case ')
						g.gen_expr(c)
						g.sb.writeln(':')
					}
				}
				g.indent++
				g.gen_stmts(branch.stmts)
				g.write_indent()
				g.sb.writeln('break;')
				g.indent--
			}
			g.write_indent()
			g.sb.writeln('}')
		}
		ast.InfixExpr {
			g.sb.write_string('(')
			g.gen_expr(node.lhs)
			op := match node.op {
				.plus { '+' }
				.minus { '-' }
				.mul { '*' }
				.div { '/' }
				.gt { '>' }
				.lt { '<' }
				.eq { '==' }
				.ne { '!=' }
				.ge { '>=' }
				.le { '<=' }
				else { '?' }
			}
			g.sb.write_string(' ${op} ')
			g.gen_expr(node.rhs)
			g.sb.write_string(')')
		}
		ast.CallExpr {
			mut name := ''
			if node.lhs is ast.Ident {
				name = node.lhs.name
			} else if node.lhs is ast.SelectorExpr {
				name = node.lhs.rhs.name
			}
			g.sb.write_string('${name}(')
			for i, arg in node.args {
				if i > 0 {
					g.sb.write_string(', ')
				}
				g.gen_expr(arg)
			}
			g.sb.write_string(')')
		}
		ast.InitExpr {
			g.sb.write_string('(${node.typ}){')
			for i, field in node.fields {
				if i > 0 {
					g.sb.write_string(', ')
				}
				g.sb.write_string('.${field.name} = ')
				g.gen_expr(field.value)
			}
			g.sb.write_string('}')
		}
		ast.SelectorExpr {
			g.gen_expr(node.lhs)
			g.sb.write_string('.')
			g.sb.write_string(node.rhs.name)
		}
		ast.IndexExpr {
			g.gen_expr(node.lhs)
			g.sb.write_string('[')
			g.gen_expr(node.expr)
			g.sb.write_string(']')
		}
		ast.PostfixExpr {
			g.gen_expr(node.expr)
			if node.op == .inc {
				g.sb.write_string('++')
			} else {
				g.sb.write_string('--')
			}
		}
		else {
			g.sb.write_string('/* expr: ${node.type_name()} */')
		}
	}
}

fn (mut g CleanCGen) write_indent() {
	for _ in 0 .. g.indent {
		g.sb.write_string('\t')
	}
}
