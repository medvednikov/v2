module veb

import fasthttp
import net.http
import time
import net
import net.urllib
import os

struct RequestParams {
	global_app         voidptr
	controllers_sorted []&ControllerPath
	routes             &map[string]Route
}

// TODO remove global hack
//__global gparams RequestParams
const gparams = RequestParams{
	routes: unsafe { nil }
}

const http_ok_response = 'HTTP/1.1 200 OK\r\nContent-Type: application/json\r\nContent-Length: 0\r\nConnection: keep-alive\r\n\r\n'.bytes()

// run_new - start a new veb server using the parallel fasthttp backend.

pub fn run_at[A, X](mut global_app A, params RunParams) ! {
	run_new[A, X](mut global_app, params.port)!
}

pub fn run_new[A, X](mut global_app A, port int) ! {
	// gapp = global_app
	if port <= 0 || port > 65535 {
		return error('invalid port number `${port}`, it should be between 1 and 65535')
	}

	// Generate routes and controllers just like the original run() function.
	routes := generate_routes[A, X](global_app)!
	controllers_sorted := check_duplicate_routes_in_controllers[A](global_app, routes)!

	unsafe {
		gparams = &RequestParams{
			global_app:         global_app
			controllers_sorted: controllers_sorted
			routes:             &routes
			// timeout_in_seconds:
		}
	}
	/*
	// This closure is the "glue". It will be executed in parallel by worker threads
	// for each incoming request.
	request_handler := fn [mut global_app, routes, controllers_sorted](req_bytes []u8, client_fd int) ![]u8 {
	}
	*/

	// Configure and run the vanilla_http_server.
	/*
	mut server := fasthttp.Server
	{
		port:            port
		request_handler: kek_handler[A, X]
	}
	*/
	mut server := fasthttp.new_server(port, parallel_request_handler[A, X]) or {
		eprintln('Failed to create server: ${err}')
		return
	}

	println('[veb] Running multi-threaded app on http://localhost:${port}/')
	flush_stdout()
	server.run() or { panic(err) }
}

// const test_text = 'test'

fn parallel_request_handler[A, X](req fasthttp.HttpRequest) ![]u8 {
	/*
	if true {
		return test_text.bytes()
	}
	*/
	// mut global_app := unsafe { &A(params.global_app) }
	//
	// mut global_app := unsafe { &A(gapp) }
	mut global_app := unsafe { &A(gparams.global_app) }
	println('parallel_request_handler() params.routes=${gparams.routes}')

	// println('global_app=$global_app')

	// println('params=$gparams')

	// println('req=$req')

	// println('buffer=${req.buffer.bytestr()}')
	s := req.buffer.bytestr()

	// method := unsafe { tos(&req.buffer[req.method.start], req.method.len) }
	// path := unsafe { tos(&req.buffer[req.path.start], req.path.len) }

	method := unsafe { tos(req.method.buf, req.method.len) }
	println('method=${method}')
	path := unsafe { tos(req.path.buf, req.path.len) }
	println('path=${path}')

	req_bytes := req.buffer
	client_fd := req.client_conn_fd

	/*

		// 1. Parse the raw request bytes into a standard `http.Request`.
		req2 := http.parse_request(req_bytes) or {
			eprintln('[veb] Failed to parse request: ${err}')
			return http_server.tiny_bad_request_response
		}
		*/

	println('s0=')
	println(s)
	println('==============')

	req2 := http.parse_request_head_str(s.clone()) or {
		eprintln('[veb] Failed to parse request: ${err}')
		println('s=')
		println(s)
		println('==============')
		return http_ok_response // http_server.tiny_bad_request_response
	}

	// println('parsed req: $req')

	// 2. Create and populate the `veb.Context`.
	completed_context := handle_request_and_route[A, X](mut global_app, req2, client_fd,
		gparams.routes, gparams.controllers_sorted)

	// 3. Serialize the final `http.Response` into a byte array.
	// Check for limitations of this synchronous backend.
	if completed_context.takeover {
		eprintln('[veb] WARNING: ctx.takeover_conn() was called, but this is not supported by this server backend. The connection will be closed after this response.')
	}

	// The vanilla_http_server expects a complete response buffer to be returned.
	println('DA RES================')
	// println(completed_context.res.body)
	return completed_context.res.bytes()

	// return  http_ok_response
}

// handle_request_and_route is a unified function that creates the context,
// runs middleware, and finds the correct route for a request.
fn handle_request_and_route[A, X](mut app A, req http.Request, client_fd int, routes &map[string]Route, controllers []&ControllerPath) &Context {
	/*
	// Create a `net.TcpConn` from the file descriptor for context compatibility.
	mut conn := &net.TcpConn{
		sock:        net.tcp_socket_from_handle_raw(client_fd)
		handle:      client_fd
		is_blocking: false // vanilla_http_server ensures this
	}
	*/

	// Create and populate the `veb.Context` from the request.
	mut url := urllib.parse(req.url) or {
		// This should be rare if http.parse_request succeeded.
		mut bad_ctx := &Context{
			req: req
			// conn: conn
		}
		bad_ctx.not_found()
		return bad_ctx
	}
	query := parse_query_from_url(url)
	form, files := parse_form_from_request(req) or {
		mut bad_ctx := &Context{
			req: req
			// conn: conn
		}
		bad_ctx.request_error('Failed to parse form data: ${err.msg()}')
		return bad_ctx
	}
	host_with_port := req.header.get(.host) or { '' }
	host, _ := urllib.split_host_port(host_with_port)

	mut ctx := &Context{
		req:            req
		page_gen_start: time.ticks()
		// conn:           conn
		query: query
		form:  form
		files: files
	}

	if connection_header := req.header.get(.connection) {
		if connection_header.to_lower() == 'close' {
			ctx.client_wants_to_close = true
		}
	}

	$if A is StaticApp {
		ctx.custom_mime_types = app.static_mime_types.clone()
	}

	// Match controller paths first
	$if A is ControllerInterface {
		if completed_context := handle_controllers[X](controllers, ctx, mut url, host) {
			return completed_context
		}
	}

	// Create a new user context and pass veb's context
	mut user_context := X{}
	user_context.Context = ctx

	println('calling handle_route')
	handle_route[A, X](mut app, mut user_context, url, host, routes)
	return &user_context.Context
}
